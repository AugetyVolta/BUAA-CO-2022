module chardet (
    input a,
    input b,
    input c
);
    
endmodule