`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:41:54 11/04/2022 
// Design Name: 
// Module Name:    ID_EX 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ID_EX(
	input 					clk,
	input						reset,
	input 					ID_EX_clr,
	input						Req,
	input       [31:0]   PC_D,
	input  		 [4:0]   A3_D,
	input 		[31:0]	RD1_D,
	input 		[31:0]	RD2_D,
	input 		 [1:0]   RD1_Sel_D,
	input			 [1:0]   RD2_Sel_D,
	input 		[31:0]	EXTImm_D,
	input			[31:0]   Instr_D,
	input			 [4:0]   A2_D,
	input 		 [4:0]	A1_D,
	input						Judge_D,
	input						BD_D,
	input			 [4:0]	Exc_Code_D,
	output reg           BD_E,
	output reg	 [4:0]	Exc_Code_E,
	output reg				Judge_E,
	output reg   [4:0]   A1_E,
	output reg   [4:0]   A2_E,
	output reg  [31:0]   Instr_E,
	output reg	[31:0] 	PC_E,
	output reg	 [4:0] 	A3_E,	//Ҫд�ļĴ�������ȥ��Ҫ���бȽ�
	output reg	[31:0] 	RD1_E,
	output reg	[31:0] 	RD2_E,
	output reg	[31:0] 	EXTImm_E,
	output reg	 [1:0] 	RD1_Sel_D_reg,
	output reg	 [1:0] 	RD2_Sel_D_reg
    );
	always@(posedge clk)begin
			if(ID_EX_clr||reset||Req)begin
				Instr_E <= 32'b0;
				PC_E <= (Req)?32'h4180:
						  (ID_EX_clr)?PC_D:
						  32'h0;//��֤���PC��ȷ
				A3_E <= 5'b0;
				RD1_E <= 32'b0;
				RD2_E <= 32'b0;
				EXTImm_E <= 32'b0;
				A2_E <= 5'b0;
				A1_E <= 5'b0;
				RD1_Sel_D_reg<= 2'b0;
				RD2_Sel_D_reg<=2'b0;
				Judge_E<=1'b0;
				BD_E<=(ID_EX_clr)?BD_D:1'b0;
				Exc_Code_E<=(ID_EX_clr)?Exc_Code_D:5'b0;
			end
			else begin
				Instr_E <= Instr_D;
				PC_E <= PC_D;
				A3_E <= A3_D;
				RD1_E <= RD1_D;
				RD2_E <= RD2_D;
				EXTImm_E <= EXTImm_D;
				A1_E <= A1_D;
				A2_E <= A2_D;
				RD1_Sel_D_reg<= RD1_Sel_D;
				RD2_Sel_D_reg<= RD2_Sel_D;
				Judge_E<=Judge_D;
				BD_E<=BD_D;
				Exc_Code_E<=Exc_Code_D;
			end
	end

endmodule
